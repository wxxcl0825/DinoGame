`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    22:04:12 12/06/2016
// Design Name:
// Module Name:    VGADEMO
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module dinosaur(input clk,
                  input [31:0]clkdiv,
                  input ena,
                  input down,
                  input jump,
                  input [11:0]lastvga_data,
                  input rstn,
                  input [8:0]row,
                  input [9:0]col,
                  output reg[11:0]vga_data,
                  output reg [9:0]x,
                  output reg [8:0]y
                 );
  wire [9:0]col_add;
  wire [8:0]row_add;
  assign col_add = 10'd72 - col + x;
  assign row_add = 9'd72 - y + row;
  reg [71:0] rom_data [0:71] = {
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000011111111111111111111111111000000,
        72'b000000000000000000000000000000000000000011111111111111111111111111000000,
        72'b000000000000000000000000000000000000000011111111111111111111111111000000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111100011111111111111111111111000,
        72'b000000000000000000000000000000000000011111100001111111111111111111111000,
        72'b000000000000000000000000000000000000011111100001111111111111111111111000,
        72'b000000000000000000000000000000000000011111100011111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111110000000000000000000,
        72'b000000000000000000000000000000000000011111111111111110000000000000000000,
        72'b000000000000000000000000000000000000011111111111111110000000000000000000,
        72'b000000000000000000000000000000000000011111111111111111111111110000000000,
        72'b000000000000000000000000000000000000011111111111111111111111111000000000,
        72'b000000000000000000000000000000000000011111111111111111111111110000000000,
        72'b000011000000000000000000000000000011111111111111100000000000000000000000,
        72'b000011100000000000000000000000000111111111111111100000000000000000000000,
        72'b000011100000000000000000000000000111111111111111100000000000000000000000,
        72'b000011100000000000000000000001111111111111111111100000000000000000000000,
        72'b000011100000000000000000000001111111111111111111100000000000000000000000,
        72'b000011100000000000000000000001111111111111111111100000000000000000000000,
        72'b000011111100000000000000111111111111111111111111111111110000000000000000,
        72'b000011111100000000000000111111111111111111111111111111110000000000000000,
        72'b000011111100000000000000111111111111111111111111111111110000000000000000,
        72'b000011111111100000001111111111111111111111111111100001110000000000000000,
        72'b000011111111100000001111111111111111111111111111100001110000000000000000,
        72'b000011111111100000001111111111111111111111111111100001110000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000000011111111111111111111111111111111111111111100000000000000000000000,
        72'b000000011111111111111111111111111111111111111100000000000000000000000000,
        72'b000000000011111111111111111111111111111111111100000000000000000000000000,
        72'b000000000001111111111111111111111111111111111100000000000000000000000000,
        72'b000000000011111111111111111111111111111111111100000000000000000000000000,
        72'b000000000000011111111111111111111111111111100000000000000000000000000000,
        72'b000000000000001111111111111111111111111111100000000000000000000000000000,
        72'b000000000000001111111111111111111111111111100000000000000000000000000000,
        72'b000000000000000001111111111111111111111100000000000000000000000000000000,
        72'b000000000000000001111111111111111111111000000000000000000000000000000000,
        72'b000000000000000001111111111111111111111000000000000000000000000000000000,
        72'b000000000000000000001111111111000111111000000000000000000000000000000000,
        72'b000000000000000000001111111111000011111000000000000000000000000000000000,
        72'b000000000000000000001111111111000111111000000000000000000000000000000000,
        72'b000000000000000000001110000000000000111000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011000000000000000000000000000000000,
        72'b000000000000000000001111111000000000011000000000000000000000000000000000,
        72'b000000000000000000001111111000000000011000000000000000000000000000000000,
        72'b000000000000000000000000000000000000011100000000000000000000000000000000,
        72'b000000000000000000000000000000000000011111100000000000000000000000000000,
        72'b000000000000000000000000000000000000011111100000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000
      };

  reg [71:0] rom2_data [0:71] = {
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000011111111111111111111111111000000,
        72'b000000000000000000000000000000000000000011111111111111111111111111000000,
        72'b000000000000000000000000000000000000000011111111111111111111111111000000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111100011111111111111111111111000,
        72'b000000000000000000000000000000000000011111100001111111111111111111111000,
        72'b000000000000000000000000000000000000011111100001111111111111111111111000,
        72'b000000000000000000000000000000000000011111100011111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111111111111111111111000,
        72'b000000000000000000000000000000000000011111111111111110000000000000000000,
        72'b000000000000000000000000000000000000011111111111111110000000000000000000,
        72'b000000000000000000000000000000000000011111111111111110000000000000000000,
        72'b000000000000000000000000000000000000011111111111111111111111110000000000,
        72'b000000000000000000000000000000000000011111111111111111111111111000000000,
        72'b000000000000000000000000000000000000011111111111111111111111110000000000,
        72'b000011000000000000000000000000000011111111111111100000000000000000000000,
        72'b000011100000000000000000000000000111111111111111100000000000000000000000,
        72'b000011100000000000000000000000000111111111111111100000000000000000000000,
        72'b000011100000000000000000000001111111111111111111100000000000000000000000,
        72'b000011100000000000000000000001111111111111111111100000000000000000000000,
        72'b000011100000000000000000000001111111111111111111100000000000000000000000,
        72'b000011111100000000000000111111111111111111111111111111110000000000000000,
        72'b000011111100000000000000111111111111111111111111111111110000000000000000,
        72'b000011111100000000000000111111111111111111111111111111110000000000000000,
        72'b000011111111100000001111111111111111111111111111100001110000000000000000,
        72'b000011111111100000001111111111111111111111111111100001110000000000000000,
        72'b000011111111100000001111111111111111111111111111100001110000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000011111111111111111111111111111111111111111111100000000000000000000000,
        72'b000000011111111111111111111111111111111111111111100000000000000000000000,
        72'b000000011111111111111111111111111111111111111100000000000000000000000000,
        72'b000000000011111111111111111111111111111111111100000000000000000000000000,
        72'b000000000001111111111111111111111111111111111100000000000000000000000000,
        72'b000000000011111111111111111111111111111111111100000000000000000000000000,
        72'b000000000000011111111111111111111111111111100000000000000000000000000000,
        72'b000000000000001111111111111111111111111111100000000000000000000000000000,
        72'b000000000000001111111111111111111111111111100000000000000000000000000000,
        72'b000000000000000001111111111111111111111100000000000000000000000000000000,
        72'b000000000000000001111111111111111111111000000000000000000000000000000000,
        72'b000000000000000001111111111111111111111000000000000000000000000000000000,
        72'b000000000000000000001111111111000111111000000000000000000000000000000000,
        72'b000000000000000000001111111111000011111000000000000000000000000000000000,
        72'b000000000000000000001111111111000111111000000000000000000000000000000000,
        72'b000000000000000000001110000000000000111000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011000000000000000000000000000000000,
        72'b000000000000000000001110000000000000011111100000000000000000000000000000,
        72'b000000000000000000001110000000000000011111100000000000000000000000000000,
        72'b000000000000000000001110000000000000000000000000000000000000000000000000,
        72'b000000000000000000001111110000000000000000000000000000000000000000000000,
        72'b000000000000000000001111110000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000
      };

  reg [71:0] down_data [0:71] = {
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000110000000000000000000000000000000000000000000000000000000000000000000,
        72'b000110000000000000000000000000000000000000000001111111111111111111000000,
        72'b000110000000000000001000000000000000000000000000111111111111111111000000,
        72'b000111111100000000001111111111111111111100000001111111111111111111000000,
        72'b000111111000000000001111111111111111111100000111111111111111111111110000,
        72'b000111111100000000001111111111111111111100000111111111111111111111111000,
        72'b000111111111111111111111111111111111111111111111100011111111111111111000,
        72'b000111111111111111111111111111111111111111111111100011111111111111111000,
        72'b000111111111111111111111111111111111111111111111100011111111111111111000,
        72'b000001111111111111111111111111111111111111111111110011111111111111111000,
        72'b000001111111111111111111111111111111111111111111111111111111111111111000,
        72'b000001111111111111111111111111111111111111111111111111111111111111111000,
        72'b000001111111111111111111111111111111111111111111111111111111111111111000,
        72'b000000011111111111111111111111111111111111111111111111111111111111111000,
        72'b000000001111111111111111111111111111111111111111111111111111111111111000,
        72'b000000001111111111111111111111111111111111111111111111111111111111111000,
        72'b000000001111111111111111111111111111111111111111111111111111111111111000,
        72'b000000000011111111111111111111111111111111111111111111111111111111111000,
        72'b000000000011111111111111111111111111111111111111111111111111111111111000,
        72'b000000000011111111111111111111111111111111111111111111111111111111111000,
        72'b000000000000111111111111111111111111111111111111111111111000000000000000,
        72'b000000000000111111111111111111111111111111111111111111111000000000000000,
        72'b000000000000111111111111111111111111111111111111111111111000000000000000,
        72'b000000000000111111111111111111111111111111111111111111111000000000000000,
        72'b000000000000000111111111111111111111111111000001111111111000000000000000,
        72'b000000000000000111111111111111111111111111000000111111111111111100000000,
        72'b000000000000000111111111111111111111111111000001111111111111111100000000,
        72'b000000000000000111111111111111111111111111000000111111111111111100000000,
        72'b000000000000000001111111111111111111111111000000000000000000000000000000,
        72'b000000000000000001111111111111111111111111000000000000000000000000000000,
        72'b000000000000000001111111111111100000001100000000000000000000000000000000,
        72'b000000000000000001111111111111100000001100000000000000000000000000000000,
        72'b000000000000000011000001111111000000001100000000000000000000000000000000,
        72'b000000000000000011000001111111000000001100000000000000000000000000000000,
        72'b000000000000000011000001111111000000001111000000000000000000000000000000,
        72'b000000000000000011000001111100000000001111000000000000000000000000000000,
        72'b000000000000000011110001111100000000001111000000000000000000000000000000,
        72'b000000000000000011110001111100000000000000000000000000000000000000000000,
        72'b000000000000000011110001111100000000000000000000000000000000000000000000,
        72'b000000000000000000000001100000000000000000000000000000000000000000000000,
        72'b000000000000000000000001100000000000000000000000000000000000000000000000,
        72'b000000000000000000000001100000000000000000000000000000000000000000000000,
        72'b000000000000000000000001100000000000000000000000000000000000000000000000,
        72'b000000000000000000000001111000000000000000000000000000000000000000000000,
        72'b000000000000000000000001111100000000000000000000000000000000000000000000,
        72'b000000000000000000000001111100000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000
      };


  reg tmp;
  reg down_flag = 1'b0;
  reg jump_flag = 1'b0;
  reg up_flag = 1'b1;
  reg [20:0]count;
  reg [7:0] cnt;
  reg [31:0] dino_count = 32'b0;
  reg dino_flag = 1'b0;
  parameter max_height = 9'd200;
  parameter min_height = 9'd329;
  parameter [8:0]state_height[0:2] = {9'd270,9'd240,9'd215};
  reg [20:0]speed = 21'd0400000;
  parameter dino_speed = 32'd040000000;
  // wire clkout;
  // Load_Gen(clk,clkdiv[17],clkdiv[18],clkout);

  always @(posedge clk or posedge rstn)
  begin
    if(rstn)
    begin
      x<=10'd41;
      y<=9'd329;
      jump_flag<=1'b0;
      down_flag<=1'b0;
      count <= 9'd0;
      dino_count <= 32'b0;
      cnt <= 0;
    end
    else
    begin
      if (!down)
      begin
        down_flag <= 1'b0;
      end
      if (down && !jump_flag)
      begin
        down_flag <= 1'b1;
      end
      if (jump && !down_flag)
      begin
        jump_flag <= 1'b1;
      end
      dino_count <= dino_count + 1;
      if(dino_count==dino_speed)
      begin
        dino_count<=0;
        dino_flag=~dino_flag;
      end
      if(jump_flag)
      begin
        count <= count + 1;
        if(y <= max_height)
        begin
          up_flag=1'b0;
        end
        if(y >= state_height[0])
        begin
          speed = 21'd0300000;
        end
        else if(y >= state_height[1])
        begin
          speed = 21'd0400000;
        end
        else if(y >= state_height[2])
        begin
          speed = 21'd0450000;
        end
		  else
		  begin
			 speed = 21'd0500000;
		  end
        if(count == speed && up_flag )
        begin
          count <= 21'd0;
          y <= y - 1;
        end
        else if(count == speed && y < min_height)
        begin
          count <=21'd0;
          y <= y + 1;
        end
        else if(count == speed)
        begin
          jump_flag <= 1'b0;
          up_flag=1'b1;
          count <= 21'd0;
        end
      end

      if(col_add < 10'd72 && row_add<9'd72 && ena)
      begin
        tmp = dino_flag?rom_data[row_add][col_add]:rom2_data[row_add][col_add];
        if(down_flag)
        begin
          tmp = down_data[row_add][col_add];
        end
        if(tmp)
        begin
          vga_data <= 12'h333;
        end
        else
        begin
          vga_data <= lastvga_data;
        end
      end
      else
      begin
        vga_data <= lastvga_data;
      end
    end
  end

endmodule
