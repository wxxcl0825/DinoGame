`timescale 1ns / 1ps
module cloud(input wire clk,
               input wire ena,
               input wire [11:0] lastvga_data,
               input wire rstn,
               input wire [8:0] row,
               input wire [9:0] col,
               input wire [20:0] speed,
               output wire [11:0] vga_data);

  parameter color = 12'hddd;
  parameter width = 78;
  parameter height = 24;


  reg [width-1:0] rom_data [0:height-1] = {
        78'b000000000000000000000000000000000000000001111111111000000000000000000000000000,
        78'b000000000000000000000000000000000111111111111111111110000000000000000000000000,
        78'b000000000000000000000000000000000111111111111111111110000000000000000000000000,
        78'b000000000000000000000000000000001111111111111111111111100000000000000000000000,
        78'b000000000000000000000000000000001111111111111001111111110000000000000000000000,
        78'b000000000000000000000000000011111111100000000000000111110000000000000000000000,
        78'b000000000000000000000000000011111111000000000000001111110000000000000000000000,
        78'b000000000000000000000000000011111111000000000000000111110000000000000000000000,
        78'b000000000000000000000000000011111110000000000000000011111111000000000000000000,
        78'b000000000000000000000000000011110000000000000000000011111111111111111000000000,
        78'b000000000000000000000000111111110000000000000000000111111111111111111000000000,
        78'b000000000000000000000000111111110000000000000000001111110111111111111000000000,
        78'b000000000000000000000111111111110000000000000000001111110111111111111111110000,
        78'b000000000011111111111111110000000000000000000000001110000000000001111111110000,
        78'b000000000011111111111111110000000000000000000000000110000000000001111111111000,
        78'b000000011111111111111111110000000000000000000000000000000000000001111111110000,
        78'b000000011111111111111111100000000000000000000000000000000000000000000001111111,
        78'b000000011111111111111111100000000000000000000000000000000000000000000001111111,
        78'b000000011111100000000000000000000000000000000000000000000000000000000001111111,
        78'b011111111110001111000000000000000000000000000000000000000000000000000001111111,
        78'b011111111111001111000000000000000000000000000000000000000000000000000000011111,
        78'b011111111111001111000000000000000000000000000000000000000000000000000000001111,
        78'b111111111111001111111111111111111111111111111111111111111111111111111111111111,
        78'b111110000000000001111111111111111111111111111111111111111111111111111111111111
      };

  reg _vga_data;

  reg [9:0] x [0:1];
  reg [8:0] y [0:1];
  reg en [0:1];

  reg [20:0] cnt;

  reg [1:0] i;
  reg [9:0] random;

  assign vga_data = (ena & _vga_data) ? color : lastvga_data;

  always @ (posedge clk or posedge rstn)
  begin
    if (rstn)
    begin
      en[0] = 0;
      en[1] = 0;
      cnt <= 0;
      x[0] = 0;
      x[1] = 320;
    end
    else
    begin
      // draw
      _vga_data = 0;
      for (i = 0; i < 2; i = i + 1)
        if (en[i] && x[i] <= col && col < x[i] + width && y[i] <= row && row < y[i] + height)
          _vga_data = _vga_data || rom_data[row - y[i]][col - x[i]];
      // emit
      if (!en[0] && random % 7 == 5)
      begin
        en[0] = 1'b1;
        x[0] = 640 + width;
        y[0] = random % 46 + 146;
        random = random * 13 + 97;
      end

      if (!en[1] && random % 5 == 1)
      begin
        en[1] = 1'b1;
        x[1] = 640 + width + random % width;
        y[1] = random % 46 + 146;
        random = random * 13 + 97;
      end

      if (cnt == speed)
      begin
        cnt <= 0;
        for (i = 0; i < 2; i = i + 1)
        begin
          if (en[i])
          begin
            x[i] = (i == 0) ? x[i] - 10'd1 : x[i] - 10'd2;
            if (x[i] == 0)
              en[i] = 0;
          end
        end
      end
      random = random * 13 + 97;
      cnt <= cnt + 1;
    end
  end

endmodule
