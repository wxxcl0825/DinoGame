module bird_cactus(
    input clk,
    input [31:0]clk_div,
    input ena,
    input [11:0] lastvga_data,
    input rstn,
    input [8:0]row,
    input [9:0]col,
    input wire [20:0] speed,
    output reg [11:0]vga_data,
    output reg crash
  );
  parameter tempvga = 12'h999;
  reg [9:0]x[0:1];
  reg [8:0]y[0:1];
  reg [9:0]col_add[0:1];
  reg [8:0]row_add[0:1];
  reg [8:0]random;
  reg [1:0]graph_type[0:1]={2'b11,2'b11};
  reg bird_flag=1'b0;

  wire [9:0]bird_width=10'd72;
  wire [8:0]bird_height=9'd49;
  wire [9:0]cactus_width=10'd56;
  wire [8:0]cactus_height=9'd56;
  wire [9:0]cactus2_width=10'd65;
  wire [8:0]cactus2_height=9'd35;

  reg [71:0] bird_data [0:48]=
      {72'b000000000000000000000000000000000000000000000000000000000000000000000000,
       72'b000000000000000000000000000000000000000000000000000000000000000000000000,
       72'b000000000000000000000000001100000000000000000000000000000000000000000000,
       72'b000000000000000000000000011100000000000000000000000000000000000000000000,
       72'b000000000000000000000000011100000000000000000000000000000000000000000000,
       72'b000000000000000000000000011110000000000000000000000000000000000000000000,
       72'b000000000000000000000000011111100000000000000000000000000000000000000000,
       72'b000000000000000000000000011111100000000000000000000000000000000000000000,
       72'b000000000000000000000000011111110000000000000000000000000000000000000000,
       72'b000000000000000000000000011111111100000000000000000000000000000000000000,
       72'b000000000000000000000000011111111100000000000000000000000000000000000000,
       72'b000000000000000000000000001111111100000000000000000000000000000000000000,
       72'b000000000000000000000000000001111110000000000000000000000000000000000000,
       72'b000000000000000011111100000001111111100000000000000000000000000000000000,
       72'b000000000000000011111100000001111111100000000000000000000000000000000000,
       72'b000000000000000011111100000001111111100000000000000000000000000000000000,
       72'b000000000000011111111100000001111111111110000000000000000000000000000000,
       72'b000000000000011111111100000001111111111100000000000000000000000000000000,
       72'b000000000000011111111100000001111111111110000000000000000000000000000000,
       72'b000000000011111111111111100001111111111111110000000000000000000000000000,
       72'b000000000011111111111111100001111111111111110000000000000000000000000000,
       72'b000000000011111111111111100001111111111111110000000000000000000000000000,
       72'b000000000111111111111111100001111111111111110000000000000000000000000000,
       72'b000000011111111111111111100001111111111111111110000000000000000000000000,
       72'b000000011111111111111111100001111111111111111110000000000000000000000000,
       72'b000000011111111111111111100001111111111111111110000000000000000000000000,
       72'b000011111111111111111111111111111111111111111110000000000000000000000000,
       72'b000011111111111111111111111111111111111111111110000000000000000000000000,
       72'b000011111111111111111111111111111111111111111110000000000000000000000000,
       72'b000000000000000000000011111111111111111111111111110000000000000000000000,
       72'b000000000000000000000011111111111111111111111111110000000000000000000000,
       72'b000000000000000000000011111111111111111111111111110000000000000000000000,
       72'b000000000000000000000000011111111111111111111111110000000000000000000000,
       72'b000000000000000000000000011111111111111111111111111111111111111111111000,
       72'b000000000000000000000000011111111111111111111111111111111111111111111000,
       72'b000000000000000000000000001111111111111111111111111111111111011111110000,
       72'b000000000000000000000000000001111111111111111111111111111110000000000000,
       72'b000000000000000000000000000001111111111111111111111111111110000000000000,
       72'b000000000000000000000000000001111111111111111111111111111110000000000000,
       72'b000000000000000000000000000000001111111111111111111111111111000000000000,
       72'b000000000000000000000000000000001111111111111111111111111111111111000000,
       72'b000000000000000000000000000000001111111111111111111111111111111110000000,
       72'b000000000000000000000000000000001111111111111111111111111111111110000000,
       72'b000000000000000000000000000000000001111111111111111111110000000000000000,
       72'b000000000000000000000000000000000001111111111111111111110000000000000000,
       72'b000000000000000000000000000000000001111111111111111111110000000000000000,
       72'b000000000000000000000000000000000000000000000000000000000000000000000000,
       72'b000000000000000000000000000000000000000000000000000000000000000000000000,
       72'b000000000000000000000000000000000000000000000000000000000000000000000000
      };
  reg [71:0] bird2_data [0:48]={
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000011111000000000000000000000000000000000000000000000000000,
        72'b000000000000000011111000000000000000000000000000000000000000000000000000,
        72'b000000000000000011111000000000000000000000000000000000000000000000000000,
        72'b000000000000001111111000000000000000000000000000000000000000000000000000,
        72'b000000000000111111111000000000000000000000000000000000000000000000000000,
        72'b000000000001111111111100000000000000000000000000000000000000000000000000,
        72'b000000000011111111111110000000000000000000000000000000000000000000000000,
        72'b000000000011111111111110000000000000000000000000000000000000000000000000,
        72'b000000000111111111111110000000000000000000000000000000000000000000000000,
        72'b000000111111111111111110000000000000000000000000000000000000000000000000,
        72'b000000111111111111111111000000000000000000000000000000000000000000000000,
        72'b000001111111111111111111110000000000000000000000000000000000000000000000,
        72'b000011111111111111111111111111111111111111111000000000000000000000000000,
        72'b000011111111111111111111111111111111111111111000000000000000000000000000,
        72'b000000000000000000000011111111111111111111111111000000000000000000000000,
        72'b000000000000000000000011111111111111111111111111000000000000000000000000,
        72'b000000000000000000000001111111111111111111111111100000000000000000000000,
        72'b000000000000000000000000011111111111111111111111100000000000000010000000,
        72'b000000000000000000000000011111111111111111111111111111111111111111000000,
        72'b000000000000000000000000000111111111111111111111111111111100000000000000,
        72'b000000000000000000000000000011111111111111111111111111111100000000000000,
        72'b000000000000000000000000000011111111111111111111111111111100000000000000,
        72'b000000000000000000000000000011111111111111111111111111111100000000000000,
        72'b000000000000000000000000000011111111111111111111111111111111111100000000,
        72'b000000000000000000000000000011111111111111111111111111111111111100000000,
        72'b000000000000000000000000000011111111111111111111111111000000000000000000,
        72'b000000000000000000000000000011111111111111111111111111000000000000000000,
        72'b000000000000000000000000000011111111111111111111111111000000000000000000,
        72'b000000000000000000000000000011111111111000000000000000000000000000000000,
        72'b000000000000000000000000000011111111111000000000000000000000000000000000,
        72'b000000000000000000000000000011111111100000000000000000000000000000000000,
        72'b000000000000000000000000000011111111100000000000000000000000000000000000,
        72'b000000000000000000000000000011111111100000000000000000000000000000000000,
        72'b000000000000000000000000000011111111000000000000000000000000000000000000,
        72'b000000000000000000000000000011111000000000000000000000000000000000000000,
        72'b000000000000000000000000000011111000000000000000000000000000000000000000,
        72'b000000000000000000000000000011111000000000000000000000000000000000000000,
        72'b000000000000000000000000000011111000000000000000000000000000000000000000,
        72'b000000000000000000000000000011111000000000000000000000000000000000000000,
        72'b000000000000000000000000000011100000000000000000000000000000000000000000,
        72'b000000000000000000000000000011000000000000000000000000000000000000000000,
        72'b000000000000000000000000000010000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000,
        72'b000000000000000000000000000000000000000000000000000000000000000000000000};
  reg [55:0] cactus_data [0:55]={
        56'b00000000000000000000000000000000000000000000000000000000,
        56'b00000000000000000000000000000000000000000000000000000000,
        56'b00000000000001110000000000000000000000011100000000000000,
        56'b00000000000011110000000000000000000000011110000000000000,
        56'b00000000001111111100000000000000000001111111100000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000100000000000001111111000000100000,
        56'b00000000000111111100001110000000000001111111000001110000,
        56'b00000000000111111100011111000000000001111111000011111000,
        56'b00000000000111111100011111000000000001111111000011110000,
        56'b00000000000111111100011111000000000001111111000011110000,
        56'b00000000000111111100011111000000000001111111000011110000,
        56'b00001000000111111100011111000001000001111111000011110000,
        56'b00001100000111111100011111000011000001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111000011110000,
        56'b00111110000111111100011111000111100001111111100011110000,
        56'b00111110000111111111111111000111100001111111111111111000,
        56'b00111110000111111111111110000111100001111111111111100000,
        56'b00111110000111111111111100000111100001111111111111100000,
        56'b00111110000111111111111000000111100001111111111110000000,
        56'b00111110000111111100000000000111100001111111100000000000,
        56'b00111110000111111100000000000111100001111111100000000000,
        56'b00111111111111111100000000000111111111111111000000000000,
        56'b00011111111111111100000000000011111111111111000000000000,
        56'b00001111111111111100000000000001111111111111000000000000,
        56'b00000111111111111100000000000000111111111111000000000000,
        56'b00000011111111111100000000000000111111111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111000000000000,
        56'b00000000000111111100000000000000000001111111100000000000,
        56'b00000000000000000000000000000000000000000000000000000000,
        56'b00000000000000000000000000000000000000000000000000000000
      };
  reg [64:0] cactus2_data [0:34]={
        65'b00000000000000000000000000000000000000000000000000000000000000000,
        65'b00000000000000000000000000000000000000000000000000000000000000000,
        65'b00000000111110000000000000000111110000000000000000011110000000000,
        65'b00000001111110000000000000000111111000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000110000111110000000000110000111111000000000,
        65'b00000001111110000110001111000111110000000000111000111111000011000,
        65'b00000001111110001111001111000111110000000000111000111111000111000,
        65'b00000001111110001110001111000111110000000000111000111111000111000,
        65'b00000001111110001110001111000111110000110000111000111111000111000,
        65'b00110001111110001110001111000111110000111000111000111111000111000,
        65'b01110001111110001110001111000111110000111000111000111111000111000,
        65'b01110001111110001110001111000111110000111000111000111111000111000,
        65'b01110001111110001110001111000111110000111000111000111111000111000,
        65'b01110001111110001110001111000111110000111000111000111111000111000,
        65'b01110001111110001110001111000111110000111000111000111111000111000,
        65'b01110001111111001111001111000111110000111000111100111111000111000,
        65'b01110001111111111100001111000111110000111000011111111111000111000,
        65'b01110001111111111000001111000111110000111000001111111111001111000,
        65'b01110001111110000000001111000111110000111000000000111111111110000,
        65'b01111001111110000000001111000111110000111000000000111111111100000,
        65'b00111111111110000000000011001111110000111000000000111111000000000,
        65'b00011111111110000000000001111111110000111000000000111111000000000,
        65'b00000001111110000000000000111111111001111000000000111111000000000,
        65'b00000001111110000000000000000111111111110000000000111111000000000,
        65'b00000001111110000000000000000111111111100000000000111111000000000,
        65'b00000001111110000000000000000111111000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000000000111110000000000000000111111000000000,
        65'b00000001111110000000000000000111111000000000000000111111000000000,
        65'b00000000000000000000000000000000000000000000000000000000000000000
      };

  reg tmp;
  reg [20:0] count;
  reg [20:0] bird_count;
  parameter bird_speed = 21'd100;

  always @(posedge clk)
  begin
      case (graph_type[0])
      2'b00:
      begin
        col_add[0] <= bird_width - col + x[0];
        row_add[0] <= bird_height - y[0] + row;
      end
      2'b01:
      begin
        col_add[0] <= bird_width - col + x[0];
        row_add[0] <= bird_height - y[0] + row;
      end
      2'b10:
      begin
        col_add[0] <= cactus_width - col + x[0];
        row_add[0] <= cactus_height + row - y[0];
      end
      2'b11:
      begin
        col_add[0] <= cactus2_width - col + x[0];
        row_add[0] <= cactus2_height + row - y[0];
      end
      default:
        ;
    endcase
    case (graph_type[1])
      2'b00:
      begin
        col_add[1] <= bird_width - col + x[1];
        row_add[1] <= bird_height - y[1] + row;
      end
      2'b01:
      begin
        col_add[1] <= bird_width - col + x[1];
        row_add[1] <= bird_height - y[1] + row;
      end
      2'b10:
      begin
        col_add[1] <= cactus_width - col + x[1];
        row_add[1] <= cactus_height + row - y[1];
      end
      2'b11:
      begin
        col_add[1] <= cactus2_width - col + x[1];
        row_add[1] <= cactus2_height + row - y[1];
      end
      default:
        ;
    endcase
    if(rstn)
    begin
      count <= 0;
      crash = 1'b0;
      x[0]<=10'd640;
      x[1]<=10'd640+10'd320;
    end
    else
    begin
      count <= count+1;

		 case(graph_type[0])
        2'b00:
        begin
          y[0]<=9'd223;
        end
        2'b01:
        begin
          y[0]<=9'd280;
        end
        2'b10:
        begin
          y[0]<=9'd331;
        end
        2'b11:
        begin
          y[0]<=9'd331;
        end
      endcase
      case(graph_type[1])
        2'b00:
        begin
          y[1]<=9'd223;
        end
        2'b01:
        begin
          y[1]<=9'd280;
        end
        2'b10:
        begin
          y[1]<=9'd331;
        end
        2'b11:
        begin
          y[1]<=9'd331;
        end
      endcase
		
      if(count==speed)
      begin
        x[0]<=x[0]-10'b1;
        x[1]<=x[1]-10'b1;
        count<=0;
        bird_count <= bird_count + 1;
      end
      if(bird_count==bird_speed)
      begin
        bird_count <= 0;
        bird_flag <= ~bird_flag;
      end

      if(x[0]==10'b0)
      begin
        x[0]<=x[0]+10'd640+random%200;
        random=random*17+47;
        graph_type[0]=random[1:0];
      end
      if(x[1]==10'b0)
      begin
        x[1]<=x[1]+10'd640+random%200;
        random=random*17+47;
        graph_type[1]=random[3:2];
      end

    end

    case (graph_type[0])
      2'b00:
      begin
        if(col_add[0] < bird_width && row_add[0] < bird_height && ena)
        begin
          tmp = bird_flag?bird_data[row_add[0]][col_add[0]]:bird2_data[row_add[0]][col_add[0]];
          if(tmp && lastvga_data==12'h333 )
          begin
            crash=1'b1;
          end
          if(tmp)
          begin
            vga_data = 12'h333;
          end
          else
          begin
            vga_data = tempvga;
          end
        end
        else
        begin
          vga_data = tempvga;
        end
      end
      2'b01:
      begin
        if(col_add[0] < bird_width && row_add[0] < bird_height && ena)
        begin
          tmp = bird_flag?bird_data[row_add[0]][col_add[0]]:bird2_data[row_add[0]][col_add[0]];
          if(tmp && lastvga_data==12'h333 )
            crash=1'b1;
          if(tmp)
          begin
            vga_data = 12'h333;
          end
          else
          begin
            vga_data = tempvga;
          end
        end
        else
        begin
          vga_data = tempvga;
        end
      end
      2'b10:
      begin
        if(col_add[0] < cactus_width && row_add[0] < cactus_height && ena)
        begin
          tmp = cactus_data[row_add[0]][col_add[0]];
          if(tmp && lastvga_data==12'h333 )
            crash=1'b1;
          if(tmp)
          begin
            vga_data = 12'h333;
          end
          else
          begin
            vga_data = tempvga;
          end
        end
        else
        begin
          vga_data = tempvga;
        end
      end
      2'b11:
      begin
        if(col_add[0] < cactus2_width && row_add[0] < cactus2_height && ena)
        begin
          tmp = cactus2_data[row_add[0]][col_add[0]];
          if(tmp && lastvga_data==12'h333 )
            crash=1'b1;
          if(tmp)
          begin
            vga_data = 12'h333;
          end
          else
          begin
            vga_data = tempvga;
          end
        end
        else
        begin
          vga_data = tempvga;
        end
      end
      default:
        ;
    endcase

    case (graph_type[1])
      2'b00:
      begin
        begin
          if(col_add[1] < bird_width && row_add[1] < bird_height && ena)
          begin
            tmp = bird_flag?bird_data[row_add[1]][col_add[1]]:bird2_data[row_add[1]][col_add[1]];
            if(tmp && lastvga_data==12'h333 )
              crash=1'b1;
            if(tmp)
            begin
              vga_data = 12'h333;
            end
          end
        end
      end
      2'b01:
      begin
        begin
          if(col_add[1] < bird_width && row_add[1] < bird_height && ena)
          begin
            tmp = bird_flag?bird_data[row_add[1]][col_add[1]]:bird2_data[row_add[1]][col_add[1]];
            if(tmp && lastvga_data==12'h333 )
              crash=1'b1;
            if(tmp)
            begin
              vga_data = 12'h333;
            end
          end
        end
      end
      2'b10:
      begin
        if(col_add[1] < cactus_width && row_add[1] < cactus_height && ena)
        begin
          tmp = cactus_data[row_add[1]][col_add[1]];
          if(tmp && lastvga_data==12'h333 )
            crash=1'b1;
          if(tmp)
          begin
            vga_data = 12'h333;
          end
        end
      end
      2'b11:
      begin
        if(col_add[1] < cactus2_width && row_add[1] < cactus2_height && ena)
        begin
          tmp = cactus2_data[row_add[1]][col_add[1]];
          if(tmp && lastvga_data==12'h333 )
            crash=1'b1;
          if(tmp)
          begin
            vga_data = 12'h333;
          end
        end
      end
      default:
        ;
    endcase
    if(vga_data==tempvga)
      vga_data=lastvga_data;
  end
endmodule
